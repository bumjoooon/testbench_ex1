class driver;
   virtual reg_if vif;
   event drv_done;
   mailbox drv_mbx;

   "
